module overlap_module_283bit(
    B2_in1,
    B2_in2,
    B2_in3,
    B2_in4,
    B2_out
    );


parameter n = 284;

input [n-2:0] B2_in1;
input [n-2:0] B2_in2;
input [n-2:0] B2_in3;
input [n-2:0] B2_in4;

output [2*n-2:0] B2_out;

assign B2_out[0] = B2_in1[0];

assign B2_out[2] = B2_in1[1]^B2_in4[0];

assign B2_out[4] = B2_in1[2]^B2_in4[1];

assign B2_out[6] = B2_in1[3]^B2_in4[2];

assign B2_out[8] = B2_in1[4]^B2_in4[3];

assign B2_out[10] = B2_in1[5]^B2_in4[4];

assign B2_out[12] = B2_in1[6]^B2_in4[5];

assign B2_out[14] = B2_in1[7]^B2_in4[6];

assign B2_out[16] = B2_in1[8]^B2_in4[7];

assign B2_out[18] = B2_in1[9]^B2_in4[8];

assign B2_out[20] = B2_in1[10]^B2_in4[9];

assign B2_out[22] = B2_in1[11]^B2_in4[10];

assign B2_out[24] = B2_in1[12]^B2_in4[11];

assign B2_out[26] = B2_in1[13]^B2_in4[12];

assign B2_out[28] = B2_in1[14]^B2_in4[13];

assign B2_out[30] = B2_in1[15]^B2_in4[14];

assign B2_out[32] = B2_in1[16]^B2_in4[15];

assign B2_out[34] = B2_in1[17]^B2_in4[16];

assign B2_out[36] = B2_in1[18]^B2_in4[17];

assign B2_out[38] = B2_in1[19]^B2_in4[18];

assign B2_out[40] = B2_in1[20]^B2_in4[19];

assign B2_out[42] = B2_in1[21]^B2_in4[20];

assign B2_out[44] = B2_in1[22]^B2_in4[21];

assign B2_out[46] = B2_in1[23]^B2_in4[22];

assign B2_out[48] = B2_in1[24]^B2_in4[23];

assign B2_out[50] = B2_in1[25]^B2_in4[24];

assign B2_out[52] = B2_in1[26]^B2_in4[25];

assign B2_out[54] = B2_in1[27]^B2_in4[26];

assign B2_out[56] = B2_in1[28]^B2_in4[27];

assign B2_out[58] = B2_in1[29]^B2_in4[28];

assign B2_out[60] = B2_in1[30]^B2_in4[29];

assign B2_out[62] = B2_in1[31]^B2_in4[30];

assign B2_out[64] = B2_in1[32]^B2_in4[31];

assign B2_out[66] = B2_in1[33]^B2_in4[32];

assign B2_out[68] = B2_in1[34]^B2_in4[33];

assign B2_out[70] = B2_in1[35]^B2_in4[34];

assign B2_out[72] = B2_in1[36]^B2_in4[35];

assign B2_out[74] = B2_in1[37]^B2_in4[36];

assign B2_out[76] = B2_in1[38]^B2_in4[37];

assign B2_out[78] = B2_in1[39]^B2_in4[38];

assign B2_out[80] = B2_in1[40]^B2_in4[39];

assign B2_out[82] = B2_in1[41]^B2_in4[40];

assign B2_out[84] = B2_in1[42]^B2_in4[41];

assign B2_out[86] = B2_in1[43]^B2_in4[42];

assign B2_out[88] = B2_in1[44]^B2_in4[43];

assign B2_out[90] = B2_in1[45]^B2_in4[44];

assign B2_out[92] = B2_in1[46]^B2_in4[45];

assign B2_out[94] = B2_in1[47]^B2_in4[46];

assign B2_out[96] = B2_in1[48]^B2_in4[47];

assign B2_out[98] = B2_in1[49]^B2_in4[48];

assign B2_out[100] = B2_in1[50]^B2_in4[49];

assign B2_out[102] = B2_in1[51]^B2_in4[50];

assign B2_out[104] = B2_in1[52]^B2_in4[51];

assign B2_out[106] = B2_in1[53]^B2_in4[52];

assign B2_out[108] = B2_in1[54]^B2_in4[53];

assign B2_out[110] = B2_in1[55]^B2_in4[54];

assign B2_out[112] = B2_in1[56]^B2_in4[55];

assign B2_out[114] = B2_in1[57]^B2_in4[56];

assign B2_out[116] = B2_in1[58]^B2_in4[57];

assign B2_out[118] = B2_in1[59]^B2_in4[58];

assign B2_out[120] = B2_in1[60]^B2_in4[59];

assign B2_out[122] = B2_in1[61]^B2_in4[60];

assign B2_out[124] = B2_in1[62]^B2_in4[61];

assign B2_out[126] = B2_in1[63]^B2_in4[62];

assign B2_out[128] = B2_in1[64]^B2_in4[63];

assign B2_out[130] = B2_in1[65]^B2_in4[64];

assign B2_out[132] = B2_in1[66]^B2_in4[65];

assign B2_out[134] = B2_in1[67]^B2_in4[66];

assign B2_out[136] = B2_in1[68]^B2_in4[67];

assign B2_out[138] = B2_in1[69]^B2_in4[68];

assign B2_out[140] = B2_in1[70]^B2_in4[69];

assign B2_out[142] = B2_in1[71]^B2_in4[70];

assign B2_out[144] = B2_in1[72]^B2_in4[71];

assign B2_out[146] = B2_in1[73]^B2_in4[72];

assign B2_out[148] = B2_in1[74]^B2_in4[73];

assign B2_out[150] = B2_in1[75]^B2_in4[74];

assign B2_out[152] = B2_in1[76]^B2_in4[75];

assign B2_out[154] = B2_in1[77]^B2_in4[76];

assign B2_out[156] = B2_in1[78]^B2_in4[77];

assign B2_out[158] = B2_in1[79]^B2_in4[78];

assign B2_out[160] = B2_in1[80]^B2_in4[79];

assign B2_out[162] = B2_in1[81]^B2_in4[80];

assign B2_out[164] = B2_in1[82]^B2_in4[81];

assign B2_out[166] = B2_in1[83]^B2_in4[82];

assign B2_out[168] = B2_in1[84]^B2_in4[83];

assign B2_out[170] = B2_in1[85]^B2_in4[84];

assign B2_out[172] = B2_in1[86]^B2_in4[85];

assign B2_out[174] = B2_in1[87]^B2_in4[86];

assign B2_out[176] = B2_in1[88]^B2_in4[87];

assign B2_out[178] = B2_in1[89]^B2_in4[88];

assign B2_out[180] = B2_in1[90]^B2_in4[89];

assign B2_out[182] = B2_in1[91]^B2_in4[90];

assign B2_out[184] = B2_in1[92]^B2_in4[91];

assign B2_out[186] = B2_in1[93]^B2_in4[92];

assign B2_out[188] = B2_in1[94]^B2_in4[93];

assign B2_out[190] = B2_in1[95]^B2_in4[94];

assign B2_out[192] = B2_in1[96]^B2_in4[95];

assign B2_out[194] = B2_in1[97]^B2_in4[96];

assign B2_out[196] = B2_in1[98]^B2_in4[97];

assign B2_out[198] = B2_in1[99]^B2_in4[98];

assign B2_out[200] = B2_in1[100]^B2_in4[99];

assign B2_out[202] = B2_in1[101]^B2_in4[100];

assign B2_out[204] = B2_in1[102]^B2_in4[101];

assign B2_out[206] = B2_in1[103]^B2_in4[102];

assign B2_out[208] = B2_in1[104]^B2_in4[103];

assign B2_out[210] = B2_in1[105]^B2_in4[104];

assign B2_out[212] = B2_in1[106]^B2_in4[105];

assign B2_out[214] = B2_in1[107]^B2_in4[106];

assign B2_out[216] = B2_in1[108]^B2_in4[107];

assign B2_out[218] = B2_in1[109]^B2_in4[108];

assign B2_out[220] = B2_in1[110]^B2_in4[109];

assign B2_out[222] = B2_in1[111]^B2_in4[110];

assign B2_out[224] = B2_in1[112]^B2_in4[111];

assign B2_out[226] = B2_in1[113]^B2_in4[112];

assign B2_out[228] = B2_in1[114]^B2_in4[113];

assign B2_out[230] = B2_in1[115]^B2_in4[114];

assign B2_out[232] = B2_in1[116]^B2_in4[115];

assign B2_out[234] = B2_in1[117]^B2_in4[116];

assign B2_out[236] = B2_in1[118]^B2_in4[117];

assign B2_out[238] = B2_in1[119]^B2_in4[118];

assign B2_out[240] = B2_in1[120]^B2_in4[119];

assign B2_out[242] = B2_in1[121]^B2_in4[120];

assign B2_out[244] = B2_in1[122]^B2_in4[121];

assign B2_out[246] = B2_in1[123]^B2_in4[122];

assign B2_out[248] = B2_in1[124]^B2_in4[123];

assign B2_out[250] = B2_in1[125]^B2_in4[124];

assign B2_out[252] = B2_in1[126]^B2_in4[125];

assign B2_out[254] = B2_in1[127]^B2_in4[126];

assign B2_out[256] = B2_in1[128]^B2_in4[127];

assign B2_out[258] = B2_in1[129]^B2_in4[128];

assign B2_out[260] = B2_in1[130]^B2_in4[129];

assign B2_out[262] = B2_in1[131]^B2_in4[130];

assign B2_out[264] = B2_in1[132]^B2_in4[131];

assign B2_out[266] = B2_in1[133]^B2_in4[132];

assign B2_out[268] = B2_in1[134]^B2_in4[133];

assign B2_out[270] = B2_in1[135]^B2_in4[134];

assign B2_out[272] = B2_in1[136]^B2_in4[135];

assign B2_out[274] = B2_in1[137]^B2_in4[136];

assign B2_out[276] = B2_in1[138]^B2_in4[137];

assign B2_out[278] = B2_in1[139]^B2_in4[138];

assign B2_out[280] = B2_in1[140]^B2_in4[139];

assign B2_out[282] = B2_in1[141]^B2_in4[140];

assign B2_out[1] = B2_in2[0]^B2_in3[0];

assign B2_out[3] = B2_in2[1]^B2_in3[1];

assign B2_out[5] = B2_in2[2]^B2_in3[2];

assign B2_out[7] = B2_in2[3]^B2_in3[3];

assign B2_out[9] = B2_in2[4]^B2_in3[4];

assign B2_out[11] = B2_in2[5]^B2_in3[5];

assign B2_out[13] = B2_in2[6]^B2_in3[6];

assign B2_out[15] = B2_in2[7]^B2_in3[7];

assign B2_out[17] = B2_in2[8]^B2_in3[8];

assign B2_out[19] = B2_in2[9]^B2_in3[9];

assign B2_out[21] = B2_in2[10]^B2_in3[10];

assign B2_out[23] = B2_in2[11]^B2_in3[11];

assign B2_out[25] = B2_in2[12]^B2_in3[12];

assign B2_out[27] = B2_in2[13]^B2_in3[13];

assign B2_out[29] = B2_in2[14]^B2_in3[14];

assign B2_out[31] = B2_in2[15]^B2_in3[15];

assign B2_out[33] = B2_in2[16]^B2_in3[16];

assign B2_out[35] = B2_in2[17]^B2_in3[17];

assign B2_out[37] = B2_in2[18]^B2_in3[18];

assign B2_out[39] = B2_in2[19]^B2_in3[19];

assign B2_out[41] = B2_in2[20]^B2_in3[20];

assign B2_out[43] = B2_in2[21]^B2_in3[21];

assign B2_out[45] = B2_in2[22]^B2_in3[22];

assign B2_out[47] = B2_in2[23]^B2_in3[23];

assign B2_out[49] = B2_in2[24]^B2_in3[24];

assign B2_out[51] = B2_in2[25]^B2_in3[25];

assign B2_out[53] = B2_in2[26]^B2_in3[26];

assign B2_out[55] = B2_in2[27]^B2_in3[27];

assign B2_out[57] = B2_in2[28]^B2_in3[28];

assign B2_out[59] = B2_in2[29]^B2_in3[29];

assign B2_out[61] = B2_in2[30]^B2_in3[30];

assign B2_out[63] = B2_in2[31]^B2_in3[31];

assign B2_out[65] = B2_in2[32]^B2_in3[32];

assign B2_out[67] = B2_in2[33]^B2_in3[33];

assign B2_out[69] = B2_in2[34]^B2_in3[34];

assign B2_out[71] = B2_in2[35]^B2_in3[35];

assign B2_out[73] = B2_in2[36]^B2_in3[36];

assign B2_out[75] = B2_in2[37]^B2_in3[37];

assign B2_out[77] = B2_in2[38]^B2_in3[38];

assign B2_out[79] = B2_in2[39]^B2_in3[39];

assign B2_out[81] = B2_in2[40]^B2_in3[40];

assign B2_out[83] = B2_in2[41]^B2_in3[41];

assign B2_out[85] = B2_in2[42]^B2_in3[42];

assign B2_out[87] = B2_in2[43]^B2_in3[43];

assign B2_out[89] = B2_in2[44]^B2_in3[44];

assign B2_out[91] = B2_in2[45]^B2_in3[45];

assign B2_out[93] = B2_in2[46]^B2_in3[46];

assign B2_out[95] = B2_in2[47]^B2_in3[47];

assign B2_out[97] = B2_in2[48]^B2_in3[48];

assign B2_out[99] = B2_in2[49]^B2_in3[49];

assign B2_out[101] = B2_in2[50]^B2_in3[50];

assign B2_out[103] = B2_in2[51]^B2_in3[51];

assign B2_out[105] = B2_in2[52]^B2_in3[52];

assign B2_out[107] = B2_in2[53]^B2_in3[53];

assign B2_out[109] = B2_in2[54]^B2_in3[54];

assign B2_out[111] = B2_in2[55]^B2_in3[55];

assign B2_out[113] = B2_in2[56]^B2_in3[56];

assign B2_out[115] = B2_in2[57]^B2_in3[57];

assign B2_out[117] = B2_in2[58]^B2_in3[58];

assign B2_out[119] = B2_in2[59]^B2_in3[59];

assign B2_out[121] = B2_in2[60]^B2_in3[60];

assign B2_out[123] = B2_in2[61]^B2_in3[61];

assign B2_out[125] = B2_in2[62]^B2_in3[62];

assign B2_out[127] = B2_in2[63]^B2_in3[63];

assign B2_out[129] = B2_in2[64]^B2_in3[64];

assign B2_out[131] = B2_in2[65]^B2_in3[65];

assign B2_out[133] = B2_in2[66]^B2_in3[66];

assign B2_out[135] = B2_in2[67]^B2_in3[67];

assign B2_out[137] = B2_in2[68]^B2_in3[68];

assign B2_out[139] = B2_in2[69]^B2_in3[69];

assign B2_out[141] = B2_in2[70]^B2_in3[70];

assign B2_out[143] = B2_in2[71]^B2_in3[71];

assign B2_out[145] = B2_in2[72]^B2_in3[72];

assign B2_out[147] = B2_in2[73]^B2_in3[73];

assign B2_out[149] = B2_in2[74]^B2_in3[74];

assign B2_out[151] = B2_in2[75]^B2_in3[75];

assign B2_out[153] = B2_in2[76]^B2_in3[76];

assign B2_out[155] = B2_in2[77]^B2_in3[77];

assign B2_out[157] = B2_in2[78]^B2_in3[78];

assign B2_out[159] = B2_in2[79]^B2_in3[79];

assign B2_out[161] = B2_in2[80]^B2_in3[80];

assign B2_out[163] = B2_in2[81]^B2_in3[81];

assign B2_out[165] = B2_in2[82]^B2_in3[82];

assign B2_out[167] = B2_in2[83]^B2_in3[83];

assign B2_out[169] = B2_in2[84]^B2_in3[84];

assign B2_out[171] = B2_in2[85]^B2_in3[85];

assign B2_out[173] = B2_in2[86]^B2_in3[86];

assign B2_out[175] = B2_in2[87]^B2_in3[87];

assign B2_out[177] = B2_in2[88]^B2_in3[88];

assign B2_out[179] = B2_in2[89]^B2_in3[89];

assign B2_out[181] = B2_in2[90]^B2_in3[90];

assign B2_out[183] = B2_in2[91]^B2_in3[91];

assign B2_out[185] = B2_in2[92]^B2_in3[92];

assign B2_out[187] = B2_in2[93]^B2_in3[93];

assign B2_out[189] = B2_in2[94]^B2_in3[94];

assign B2_out[191] = B2_in2[95]^B2_in3[95];

assign B2_out[193] = B2_in2[96]^B2_in3[96];

assign B2_out[195] = B2_in2[97]^B2_in3[97];

assign B2_out[197] = B2_in2[98]^B2_in3[98];

assign B2_out[199] = B2_in2[99]^B2_in3[99];

assign B2_out[201] = B2_in2[100]^B2_in3[100];

assign B2_out[203] = B2_in2[101]^B2_in3[101];

assign B2_out[205] = B2_in2[102]^B2_in3[102];

assign B2_out[207] = B2_in2[103]^B2_in3[103];

assign B2_out[209] = B2_in2[104]^B2_in3[104];

assign B2_out[211] = B2_in2[105]^B2_in3[105];

assign B2_out[213] = B2_in2[106]^B2_in3[106];

assign B2_out[215] = B2_in2[107]^B2_in3[107];

assign B2_out[217] = B2_in2[108]^B2_in3[108];

assign B2_out[219] = B2_in2[109]^B2_in3[109];

assign B2_out[221] = B2_in2[110]^B2_in3[110];

assign B2_out[223] = B2_in2[111]^B2_in3[111];

assign B2_out[225] = B2_in2[112]^B2_in3[112];

assign B2_out[227] = B2_in2[113]^B2_in3[113];

assign B2_out[229] = B2_in2[114]^B2_in3[114];

assign B2_out[231] = B2_in2[115]^B2_in3[115];

assign B2_out[233] = B2_in2[116]^B2_in3[116];

assign B2_out[235] = B2_in2[117]^B2_in3[117];

assign B2_out[237] = B2_in2[118]^B2_in3[118];

assign B2_out[239] = B2_in2[119]^B2_in3[119];

assign B2_out[241] = B2_in2[120]^B2_in3[120];

assign B2_out[243] = B2_in2[121]^B2_in3[121];

assign B2_out[245] = B2_in2[122]^B2_in3[122];

assign B2_out[247] = B2_in2[123]^B2_in3[123];

assign B2_out[249] = B2_in2[124]^B2_in3[124];

assign B2_out[251] = B2_in2[125]^B2_in3[125];

assign B2_out[253] = B2_in2[126]^B2_in3[126];

assign B2_out[255] = B2_in2[127]^B2_in3[127];

assign B2_out[257] = B2_in2[128]^B2_in3[128];

assign B2_out[259] = B2_in2[129]^B2_in3[129];

assign B2_out[261] = B2_in2[130]^B2_in3[130];

assign B2_out[263] = B2_in2[131]^B2_in3[131];

assign B2_out[265] = B2_in2[132]^B2_in3[132];

assign B2_out[267] = B2_in2[133]^B2_in3[133];

assign B2_out[269] = B2_in2[134]^B2_in3[134];

assign B2_out[271] = B2_in2[135]^B2_in3[135];

assign B2_out[273] = B2_in2[136]^B2_in3[136];

assign B2_out[275] = B2_in2[137]^B2_in3[137];

assign B2_out[277] = B2_in2[138]^B2_in3[138];

assign B2_out[279] = B2_in2[139]^B2_in3[139];

assign B2_out[281] = B2_in2[140]^B2_in3[140];

assign B2_out[283] = B2_in2[141]^B2_in3[141];

assign B2_out[285] = B2_in2[142]^B2_in3[142];

assign B2_out[287] = B2_in2[143]^B2_in3[143];

assign B2_out[289] = B2_in2[144]^B2_in3[144];

assign B2_out[291] = B2_in2[145]^B2_in3[145];

assign B2_out[293] = B2_in2[146]^B2_in3[146];

assign B2_out[295] = B2_in2[147]^B2_in3[147];

assign B2_out[297] = B2_in2[148]^B2_in3[148];

assign B2_out[299] = B2_in2[149]^B2_in3[149];

assign B2_out[301] = B2_in2[150]^B2_in3[150];

assign B2_out[303] = B2_in2[151]^B2_in3[151];

assign B2_out[305] = B2_in2[152]^B2_in3[152];

assign B2_out[307] = B2_in2[153]^B2_in3[153];

assign B2_out[309] = B2_in2[154]^B2_in3[154];

assign B2_out[311] = B2_in2[155]^B2_in3[155];

assign B2_out[313] = B2_in2[156]^B2_in3[156];

assign B2_out[315] = B2_in2[157]^B2_in3[157];

assign B2_out[317] = B2_in2[158]^B2_in3[158];

assign B2_out[319] = B2_in2[159]^B2_in3[159];

assign B2_out[321] = B2_in2[160]^B2_in3[160];

assign B2_out[323] = B2_in2[161]^B2_in3[161];

assign B2_out[325] = B2_in2[162]^B2_in3[162];

assign B2_out[327] = B2_in2[163]^B2_in3[163];

assign B2_out[329] = B2_in2[164]^B2_in3[164];

assign B2_out[331] = B2_in2[165]^B2_in3[165];

assign B2_out[333] = B2_in2[166]^B2_in3[166];

assign B2_out[335] = B2_in2[167]^B2_in3[167];

assign B2_out[337] = B2_in2[168]^B2_in3[168];

assign B2_out[339] = B2_in2[169]^B2_in3[169];

assign B2_out[341] = B2_in2[170]^B2_in3[170];

assign B2_out[343] = B2_in2[171]^B2_in3[171];

assign B2_out[345] = B2_in2[172]^B2_in3[172];

assign B2_out[347] = B2_in2[173]^B2_in3[173];

assign B2_out[349] = B2_in2[174]^B2_in3[174];

assign B2_out[351] = B2_in2[175]^B2_in3[175];

assign B2_out[353] = B2_in2[176]^B2_in3[176];

assign B2_out[355] = B2_in2[177]^B2_in3[177];

assign B2_out[357] = B2_in2[178]^B2_in3[178];

assign B2_out[359] = B2_in2[179]^B2_in3[179];

assign B2_out[361] = B2_in2[180]^B2_in3[180];

assign B2_out[363] = B2_in2[181]^B2_in3[181];

assign B2_out[365] = B2_in2[182]^B2_in3[182];

assign B2_out[367] = B2_in2[183]^B2_in3[183];

assign B2_out[369] = B2_in2[184]^B2_in3[184];

assign B2_out[371] = B2_in2[185]^B2_in3[185];

assign B2_out[373] = B2_in2[186]^B2_in3[186];

assign B2_out[375] = B2_in2[187]^B2_in3[187];

assign B2_out[377] = B2_in2[188]^B2_in3[188];

assign B2_out[379] = B2_in2[189]^B2_in3[189];

assign B2_out[381] = B2_in2[190]^B2_in3[190];

assign B2_out[383] = B2_in2[191]^B2_in3[191];

assign B2_out[385] = B2_in2[192]^B2_in3[192];

assign B2_out[387] = B2_in2[193]^B2_in3[193];

assign B2_out[389] = B2_in2[194]^B2_in3[194];

assign B2_out[391] = B2_in2[195]^B2_in3[195];

assign B2_out[393] = B2_in2[196]^B2_in3[196];

assign B2_out[395] = B2_in2[197]^B2_in3[197];

assign B2_out[397] = B2_in2[198]^B2_in3[198];

assign B2_out[399] = B2_in2[199]^B2_in3[199];

assign B2_out[401] = B2_in2[200]^B2_in3[200];

assign B2_out[403] = B2_in2[201]^B2_in3[201];

assign B2_out[405] = B2_in2[202]^B2_in3[202];

assign B2_out[407] = B2_in2[203]^B2_in3[203];

assign B2_out[409] = B2_in2[204]^B2_in3[204];

assign B2_out[411] = B2_in2[205]^B2_in3[205];

assign B2_out[413] = B2_in2[206]^B2_in3[206];

assign B2_out[415] = B2_in2[207]^B2_in3[207];

assign B2_out[417] = B2_in2[208]^B2_in3[208];

assign B2_out[419] = B2_in2[209]^B2_in3[209];

assign B2_out[421] = B2_in2[210]^B2_in3[210];

assign B2_out[423] = B2_in2[211]^B2_in3[211];

assign B2_out[425] = B2_in2[212]^B2_in3[212];

assign B2_out[427] = B2_in2[213]^B2_in3[213];

assign B2_out[429] = B2_in2[214]^B2_in3[214];

assign B2_out[431] = B2_in2[215]^B2_in3[215];

assign B2_out[433] = B2_in2[216]^B2_in3[216];

assign B2_out[435] = B2_in2[217]^B2_in3[217];

assign B2_out[437] = B2_in2[218]^B2_in3[218];

assign B2_out[439] = B2_in2[219]^B2_in3[219];

assign B2_out[441] = B2_in2[220]^B2_in3[220];

assign B2_out[443] = B2_in2[221]^B2_in3[221];

assign B2_out[445] = B2_in2[222]^B2_in3[222];

assign B2_out[447] = B2_in2[223]^B2_in3[223];

assign B2_out[449] = B2_in2[224]^B2_in3[224];

assign B2_out[451] = B2_in2[225]^B2_in3[225];

assign B2_out[453] = B2_in2[226]^B2_in3[226];

assign B2_out[455] = B2_in2[227]^B2_in3[227];

assign B2_out[457] = B2_in2[228]^B2_in3[228];

assign B2_out[459] = B2_in2[229]^B2_in3[229];

assign B2_out[461] = B2_in2[230]^B2_in3[230];

assign B2_out[463] = B2_in2[231]^B2_in3[231];

assign B2_out[465] = B2_in2[232]^B2_in3[232];

assign B2_out[467] = B2_in2[233]^B2_in3[233];

assign B2_out[469] = B2_in2[234]^B2_in3[234];

assign B2_out[471] = B2_in2[235]^B2_in3[235];

assign B2_out[473] = B2_in2[236]^B2_in3[236];

assign B2_out[475] = B2_in2[237]^B2_in3[237];

assign B2_out[477] = B2_in2[238]^B2_in3[238];

assign B2_out[479] = B2_in2[239]^B2_in3[239];

assign B2_out[481] = B2_in2[240]^B2_in3[240];

assign B2_out[483] = B2_in2[241]^B2_in3[241];

assign B2_out[485] = B2_in2[242]^B2_in3[242];

assign B2_out[487] = B2_in2[243]^B2_in3[243];

assign B2_out[489] = B2_in2[244]^B2_in3[244];

assign B2_out[491] = B2_in2[245]^B2_in3[245];

assign B2_out[493] = B2_in2[246]^B2_in3[246];

assign B2_out[495] = B2_in2[247]^B2_in3[247];

assign B2_out[497] = B2_in2[248]^B2_in3[248];

assign B2_out[499] = B2_in2[249]^B2_in3[249];

assign B2_out[501] = B2_in2[250]^B2_in3[250];

assign B2_out[503] = B2_in2[251]^B2_in3[251];

assign B2_out[505] = B2_in2[252]^B2_in3[252];

assign B2_out[507] = B2_in2[253]^B2_in3[253];

assign B2_out[509] = B2_in2[254]^B2_in3[254];

assign B2_out[511] = B2_in2[255]^B2_in3[255];

assign B2_out[513] = B2_in2[256]^B2_in3[256];

assign B2_out[515] = B2_in2[257]^B2_in3[257];

assign B2_out[517] = B2_in2[258]^B2_in3[258];

assign B2_out[519] = B2_in2[259]^B2_in3[259];

assign B2_out[521] = B2_in2[260]^B2_in3[260];

assign B2_out[523] = B2_in2[261]^B2_in3[261];

assign B2_out[525] = B2_in2[262]^B2_in3[262];

assign B2_out[527] = B2_in2[263]^B2_in3[263];

assign B2_out[529] = B2_in2[264]^B2_in3[264];

assign B2_out[531] = B2_in2[265]^B2_in3[265];

assign B2_out[533] = B2_in2[266]^B2_in3[266];

assign B2_out[535] = B2_in2[267]^B2_in3[267];

assign B2_out[537] = B2_in2[268]^B2_in3[268];

assign B2_out[539] = B2_in2[269]^B2_in3[269];

assign B2_out[541] = B2_in2[270]^B2_in3[270];

assign B2_out[543] = B2_in2[271]^B2_in3[271];

assign B2_out[545] = B2_in2[272]^B2_in3[272];

assign B2_out[547] = B2_in2[273]^B2_in3[273];

assign B2_out[549] = B2_in2[274]^B2_in3[274];

assign B2_out[551] = B2_in2[275]^B2_in3[275];

assign B2_out[553] = B2_in2[276]^B2_in3[276];

assign B2_out[555] = B2_in2[277]^B2_in3[277];

assign B2_out[557] = B2_in2[278]^B2_in3[278];

assign B2_out[559] = B2_in2[279]^B2_in3[279];

assign B2_out[561] = B2_in2[280]^B2_in3[280];

assign B2_out[563] = B2_in2[281]^B2_in3[281];

assign B2_out[565] = B2_in2[282]^B2_in3[282];

assign B2_out[284] = B2_in1[142]^B2_in4[141];

assign B2_out[286] = B2_in1[143]^B2_in4[142];

assign B2_out[288] = B2_in1[144]^B2_in4[143];

assign B2_out[290] = B2_in1[145]^B2_in4[144];

assign B2_out[292] = B2_in1[146]^B2_in4[145];

assign B2_out[294] = B2_in1[147]^B2_in4[146];

assign B2_out[296] = B2_in1[148]^B2_in4[147];

assign B2_out[298] = B2_in1[149]^B2_in4[148];

assign B2_out[300] = B2_in1[150]^B2_in4[149];

assign B2_out[302] = B2_in1[151]^B2_in4[150];

assign B2_out[304] = B2_in1[152]^B2_in4[151];

assign B2_out[306] = B2_in1[153]^B2_in4[152];

assign B2_out[308] = B2_in1[154]^B2_in4[153];

assign B2_out[310] = B2_in1[155]^B2_in4[154];

assign B2_out[312] = B2_in1[156]^B2_in4[155];

assign B2_out[314] = B2_in1[157]^B2_in4[156];

assign B2_out[316] = B2_in1[158]^B2_in4[157];

assign B2_out[318] = B2_in1[159]^B2_in4[158];

assign B2_out[320] = B2_in1[160]^B2_in4[159];

assign B2_out[322] = B2_in1[161]^B2_in4[160];

assign B2_out[324] = B2_in1[162]^B2_in4[161];

assign B2_out[326] = B2_in1[163]^B2_in4[162];

assign B2_out[328] = B2_in1[164]^B2_in4[163];

assign B2_out[330] = B2_in1[165]^B2_in4[164];

assign B2_out[332] = B2_in1[166]^B2_in4[165];

assign B2_out[334] = B2_in1[167]^B2_in4[166];

assign B2_out[336] = B2_in1[168]^B2_in4[167];

assign B2_out[338] = B2_in1[169]^B2_in4[168];

assign B2_out[340] = B2_in1[170]^B2_in4[169];

assign B2_out[342] = B2_in1[171]^B2_in4[170];

assign B2_out[344] = B2_in1[172]^B2_in4[171];

assign B2_out[346] = B2_in1[173]^B2_in4[172];

assign B2_out[348] = B2_in1[174]^B2_in4[173];

assign B2_out[350] = B2_in1[175]^B2_in4[174];

assign B2_out[352] = B2_in1[176]^B2_in4[175];

assign B2_out[354] = B2_in1[177]^B2_in4[176];

assign B2_out[356] = B2_in1[178]^B2_in4[177];

assign B2_out[358] = B2_in1[179]^B2_in4[178];

assign B2_out[360] = B2_in1[180]^B2_in4[179];

assign B2_out[362] = B2_in1[181]^B2_in4[180];

assign B2_out[364] = B2_in1[182]^B2_in4[181];

assign B2_out[366] = B2_in1[183]^B2_in4[182];

assign B2_out[368] = B2_in1[184]^B2_in4[183];

assign B2_out[370] = B2_in1[185]^B2_in4[184];

assign B2_out[372] = B2_in1[186]^B2_in4[185];

assign B2_out[374] = B2_in1[187]^B2_in4[186];

assign B2_out[376] = B2_in1[188]^B2_in4[187];

assign B2_out[378] = B2_in1[189]^B2_in4[188];

assign B2_out[380] = B2_in1[190]^B2_in4[189];

assign B2_out[382] = B2_in1[191]^B2_in4[190];

assign B2_out[384] = B2_in1[192]^B2_in4[191];

assign B2_out[386] = B2_in1[193]^B2_in4[192];

assign B2_out[388] = B2_in1[194]^B2_in4[193];

assign B2_out[390] = B2_in1[195]^B2_in4[194];

assign B2_out[392] = B2_in1[196]^B2_in4[195];

assign B2_out[394] = B2_in1[197]^B2_in4[196];

assign B2_out[396] = B2_in1[198]^B2_in4[197];

assign B2_out[398] = B2_in1[199]^B2_in4[198];

assign B2_out[400] = B2_in1[200]^B2_in4[199];

assign B2_out[402] = B2_in1[201]^B2_in4[200];

assign B2_out[404] = B2_in1[202]^B2_in4[201];

assign B2_out[406] = B2_in1[203]^B2_in4[202];

assign B2_out[408] = B2_in1[204]^B2_in4[203];

assign B2_out[410] = B2_in1[205]^B2_in4[204];

assign B2_out[412] = B2_in1[206]^B2_in4[205];

assign B2_out[414] = B2_in1[207]^B2_in4[206];

assign B2_out[416] = B2_in1[208]^B2_in4[207];

assign B2_out[418] = B2_in1[209]^B2_in4[208];

assign B2_out[420] = B2_in1[210]^B2_in4[209];

assign B2_out[422] = B2_in1[211]^B2_in4[210];

assign B2_out[424] = B2_in1[212]^B2_in4[211];

assign B2_out[426] = B2_in1[213]^B2_in4[212];

assign B2_out[428] = B2_in1[214]^B2_in4[213];

assign B2_out[430] = B2_in1[215]^B2_in4[214];

assign B2_out[432] = B2_in1[216]^B2_in4[215];

assign B2_out[434] = B2_in1[217]^B2_in4[216];

assign B2_out[436] = B2_in1[218]^B2_in4[217];

assign B2_out[438] = B2_in1[219]^B2_in4[218];

assign B2_out[440] = B2_in1[220]^B2_in4[219];

assign B2_out[442] = B2_in1[221]^B2_in4[220];

assign B2_out[444] = B2_in1[222]^B2_in4[221];

assign B2_out[446] = B2_in1[223]^B2_in4[222];

assign B2_out[448] = B2_in1[224]^B2_in4[223];

assign B2_out[450] = B2_in1[225]^B2_in4[224];

assign B2_out[452] = B2_in1[226]^B2_in4[225];

assign B2_out[454] = B2_in1[227]^B2_in4[226];

assign B2_out[456] = B2_in1[228]^B2_in4[227];

assign B2_out[458] = B2_in1[229]^B2_in4[228];

assign B2_out[460] = B2_in1[230]^B2_in4[229];

assign B2_out[462] = B2_in1[231]^B2_in4[230];

assign B2_out[464] = B2_in1[232]^B2_in4[231];

assign B2_out[466] = B2_in1[233]^B2_in4[232];

assign B2_out[468] = B2_in1[234]^B2_in4[233];

assign B2_out[470] = B2_in1[235]^B2_in4[234];

assign B2_out[472] = B2_in1[236]^B2_in4[235];

assign B2_out[474] = B2_in1[237]^B2_in4[236];

assign B2_out[476] = B2_in1[238]^B2_in4[237];

assign B2_out[478] = B2_in1[239]^B2_in4[238];

assign B2_out[480] = B2_in1[240]^B2_in4[239];

assign B2_out[482] = B2_in1[241]^B2_in4[240];

assign B2_out[484] = B2_in1[242]^B2_in4[241];

assign B2_out[486] = B2_in1[243]^B2_in4[242];

assign B2_out[488] = B2_in1[244]^B2_in4[243];

assign B2_out[490] = B2_in1[245]^B2_in4[244];

assign B2_out[492] = B2_in1[246]^B2_in4[245];

assign B2_out[494] = B2_in1[247]^B2_in4[246];

assign B2_out[496] = B2_in1[248]^B2_in4[247];

assign B2_out[498] = B2_in1[249]^B2_in4[248];

assign B2_out[500] = B2_in1[250]^B2_in4[249];

assign B2_out[502] = B2_in1[251]^B2_in4[250];

assign B2_out[504] = B2_in1[252]^B2_in4[251];

assign B2_out[506] = B2_in1[253]^B2_in4[252];

assign B2_out[508] = B2_in1[254]^B2_in4[253];

assign B2_out[510] = B2_in1[255]^B2_in4[254];

assign B2_out[512] = B2_in1[256]^B2_in4[255];

assign B2_out[514] = B2_in1[257]^B2_in4[256];

assign B2_out[516] = B2_in1[258]^B2_in4[257];

assign B2_out[518] = B2_in1[259]^B2_in4[258];

assign B2_out[520] = B2_in1[260]^B2_in4[259];

assign B2_out[522] = B2_in1[261]^B2_in4[260];

assign B2_out[524] = B2_in1[262]^B2_in4[261];

assign B2_out[526] = B2_in1[263]^B2_in4[262];

assign B2_out[528] = B2_in1[264]^B2_in4[263];

assign B2_out[530] = B2_in1[265]^B2_in4[264];

assign B2_out[532] = B2_in1[266]^B2_in4[265];

assign B2_out[534] = B2_in1[267]^B2_in4[266];

assign B2_out[536] = B2_in1[268]^B2_in4[267];

assign B2_out[538] = B2_in1[269]^B2_in4[268];

assign B2_out[540] = B2_in1[270]^B2_in4[269];

assign B2_out[542] = B2_in1[271]^B2_in4[270];

assign B2_out[544] = B2_in1[272]^B2_in4[271];

assign B2_out[546] = B2_in1[273]^B2_in4[272];

assign B2_out[548] = B2_in1[274]^B2_in4[273];

assign B2_out[550] = B2_in1[275]^B2_in4[274];

assign B2_out[552] = B2_in1[276]^B2_in4[275];

assign B2_out[554] = B2_in1[277]^B2_in4[276];

assign B2_out[556] = B2_in1[278]^B2_in4[277];

assign B2_out[558] = B2_in1[279]^B2_in4[278];

assign B2_out[560] = B2_in1[280]^B2_in4[279];

assign B2_out[562] = B2_in1[281]^B2_in4[280];

assign B2_out[564] = B2_in1[282]^B2_in4[281];

assign B2_out[566] = B2_in4[282];

endmodule